class interface;
  logic [7:0] a;
  logic [7:0] b;
  logic [7:0] y;
endinterface
