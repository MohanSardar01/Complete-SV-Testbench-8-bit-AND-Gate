module andt (
  input [7:0] a,b;
  outpur [7:0] y
);
  
  assign y = a & b;
  
endmodule
