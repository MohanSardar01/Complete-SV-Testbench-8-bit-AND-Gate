class environment;
  
endclass
